* Spice netlister for gnetlist
R1 N001 0 1k
R2 Vout N001 4k
R3 N003 N002 250
R 0 N003 250
C1 N002 0 1m
C2 Vout N003 1m
XU1 N002 N001 Vcc -Vcc Vout LM741/NS
V1 Vcc 0 12
V2 0 -Vcc 12
.PRINT TRAN t V(vout)
.tran 0.02ms 25s
.include LM741.MOD
*.backanno
*.control
*run
*plot V(vout)
*.endc
.end
